* Simple RC test for Xyce
V1 in 0 AC 1
R1 in out 1k
C1 out 0 1u

.ac dec 10 10 1e6
.print ac V(out)
.end
